* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__schmittbuf_1 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
rI39 net069 VGND sky130_fd_pr__res_generic_nd__hv m=1 w=0.29 l=1.355 isHV=TRUE
rI38 VPWR net32 sky130_fd_pr__res_generic_pd__hv m=1 w=0.29 l=3.11 isHV=TRUE
MI5 net32 net36 net40 VNB nfet_g5v0d10v5 m=1 w=0.42 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 net36 A net40 VNB nfet_g5v0d10v5 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 net40 A VGND VNB nfet_g5v0d10v5 m=1 w=0.42 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X net36 VGND VNB nfet_g5v0d10v5 m=1 w=0.75 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI6 net069 net36 net56 VPB pfet_g5v0d10v5 m=1 w=0.75 l=0.5 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP0 VPWR A net56 VPB pfet_g5v0d10v5 m=1 w=0.75 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 net56 A net36 VPB pfet_g5v0d10v5 m=1 w=0.75 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X net36 VPWR VPB pfet_g5v0d10v5 m=1 w=1.5 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_hvl__schmittbuf_1
