/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1_PP_BLACKBOX_V
`define SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1_PP_BLACKBOX_V

/**
 * lsbufhv2hv_hl: Level shifting buffer, High Voltage to High Voltage,
 *                Higher Voltage to Lower Voltage.
 *
 * Verilog stub definition (black box with power pins).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_sc_hvl__lsbufhv2hv_hl_1 (
    X       ,
    A       ,
    VPWR    ,
    VGND    ,
    LOWHVPWR,
    VPB     ,
    VNB
);

    output X       ;
    input  A       ;
    input  VPWR    ;
    input  VGND    ;
    input  LOWHVPWR;
    input  VPB     ;
    input  VNB     ;
endmodule

`default_nettype wire
`endif  // SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1_PP_BLACKBOX_V
